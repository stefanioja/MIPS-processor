module AND(Input1,
           Input2,
           Output);
  
  input Input1;
  input Input2;
  output Output;
  
  assign Output = Input1 & Input2;
endmodule